// compression.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module compression (
		input  wire        clk_clk,          //       clk.clk
		output wire [7:0]  leds_w_export,    //    leds_w.export
		input  wire [31:0] line1_1_in_port,  //   line1_1.in_port
		output wire [31:0] line1_1_out_port, //          .out_port
		input  wire [31:0] line1_2_in_port,  //   line1_2.in_port
		output wire [31:0] line1_2_out_port, //          .out_port
		input  wire [31:0] line2_1_in_port,  //   line2_1.in_port
		output wire [31:0] line2_1_out_port, //          .out_port
		input  wire [31:0] line2_2_in_port,  //   line2_2.in_port
		output wire [31:0] line2_2_out_port, //          .out_port
		input  wire [31:0] line3_1_in_port,  //   line3_1.in_port
		output wire [31:0] line3_1_out_port, //          .out_port
		input  wire [31:0] line3_2_in_port,  //   line3_2.in_port
		output wire [31:0] line3_2_out_port, //          .out_port
		input  wire [31:0] line4_1_in_port,  //   line4_1.in_port
		output wire [31:0] line4_1_out_port, //          .out_port
		input  wire [31:0] line4_2_in_port,  //   line4_2.in_port
		output wire [31:0] line4_2_out_port, //          .out_port
		input  wire [31:0] line5_1_in_port,  //   line5_1.in_port
		output wire [31:0] line5_1_out_port, //          .out_port
		input  wire [31:0] line5_2_in_port,  //   line5_2.in_port
		output wire [31:0] line5_2_out_port, //          .out_port
		input  wire [31:0] line6_1_in_port,  //   line6_1.in_port
		output wire [31:0] line6_1_out_port, //          .out_port
		input  wire [31:0] line6_2_in_port,  //   line6_2.in_port
		output wire [31:0] line6_2_out_port, //          .out_port
		input  wire [31:0] line7_1_in_port,  //   line7_1.in_port
		output wire [31:0] line7_1_out_port, //          .out_port
		input  wire [31:0] line7_2_in_port,  //   line7_2.in_port
		output wire [31:0] line7_2_out_port, //          .out_port
		input  wire [31:0] line8_1_in_port,  //   line8_1.in_port
		output wire [31:0] line8_1_out_port, //          .out_port
		input  wire [31:0] line8_2_in_port,  //   line8_2.in_port
		output wire [31:0] line8_2_out_port, //          .out_port
		input  wire        reset_reset_n,    //     reset.reset_n
		output wire [11:0] sdram_addr,       //     sdram.addr
		output wire [1:0]  sdram_ba,         //          .ba
		output wire        sdram_cas_n,      //          .cas_n
		output wire        sdram_cke,        //          .cke
		output wire        sdram_cs_n,       //          .cs_n
		inout  wire [31:0] sdram_dq,         //          .dq
		output wire [3:0]  sdram_dqm,        //          .dqm
		output wire        sdram_ras_n,      //          .ras_n
		output wire        sdram_we_n,       //          .we_n
		output wire        sdram_pll_clk     // sdram_pll.clk
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;             // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;              // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                 // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;            // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                      // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                        // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                         // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                           // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                       // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;          // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;            // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;         // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_controller_s1_address;             // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;          // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;       // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;               // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;           // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;          // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;            // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;             // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;          // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;               // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;           // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;               // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_line1_1_s1_chipselect;                   // mm_interconnect_0:Line1_1_s1_chipselect -> Line1_1:chipselect
	wire  [31:0] mm_interconnect_0_line1_1_s1_readdata;                     // Line1_1:readdata -> mm_interconnect_0:Line1_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line1_1_s1_address;                      // mm_interconnect_0:Line1_1_s1_address -> Line1_1:address
	wire         mm_interconnect_0_line1_1_s1_write;                        // mm_interconnect_0:Line1_1_s1_write -> Line1_1:write_n
	wire  [31:0] mm_interconnect_0_line1_1_s1_writedata;                    // mm_interconnect_0:Line1_1_s1_writedata -> Line1_1:writedata
	wire         mm_interconnect_0_line1_2_s1_chipselect;                   // mm_interconnect_0:Line1_2_s1_chipselect -> Line1_2:chipselect
	wire  [31:0] mm_interconnect_0_line1_2_s1_readdata;                     // Line1_2:readdata -> mm_interconnect_0:Line1_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line1_2_s1_address;                      // mm_interconnect_0:Line1_2_s1_address -> Line1_2:address
	wire         mm_interconnect_0_line1_2_s1_write;                        // mm_interconnect_0:Line1_2_s1_write -> Line1_2:write_n
	wire  [31:0] mm_interconnect_0_line1_2_s1_writedata;                    // mm_interconnect_0:Line1_2_s1_writedata -> Line1_2:writedata
	wire         mm_interconnect_0_line8_2_s1_chipselect;                   // mm_interconnect_0:Line8_2_s1_chipselect -> Line8_2:chipselect
	wire  [31:0] mm_interconnect_0_line8_2_s1_readdata;                     // Line8_2:readdata -> mm_interconnect_0:Line8_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line8_2_s1_address;                      // mm_interconnect_0:Line8_2_s1_address -> Line8_2:address
	wire         mm_interconnect_0_line8_2_s1_write;                        // mm_interconnect_0:Line8_2_s1_write -> Line8_2:write_n
	wire  [31:0] mm_interconnect_0_line8_2_s1_writedata;                    // mm_interconnect_0:Line8_2_s1_writedata -> Line8_2:writedata
	wire         mm_interconnect_0_line8_1_s1_chipselect;                   // mm_interconnect_0:Line8_1_s1_chipselect -> Line8_1:chipselect
	wire  [31:0] mm_interconnect_0_line8_1_s1_readdata;                     // Line8_1:readdata -> mm_interconnect_0:Line8_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line8_1_s1_address;                      // mm_interconnect_0:Line8_1_s1_address -> Line8_1:address
	wire         mm_interconnect_0_line8_1_s1_write;                        // mm_interconnect_0:Line8_1_s1_write -> Line8_1:write_n
	wire  [31:0] mm_interconnect_0_line8_1_s1_writedata;                    // mm_interconnect_0:Line8_1_s1_writedata -> Line8_1:writedata
	wire         mm_interconnect_0_line7_2_s1_chipselect;                   // mm_interconnect_0:Line7_2_s1_chipselect -> Line7_2:chipselect
	wire  [31:0] mm_interconnect_0_line7_2_s1_readdata;                     // Line7_2:readdata -> mm_interconnect_0:Line7_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line7_2_s1_address;                      // mm_interconnect_0:Line7_2_s1_address -> Line7_2:address
	wire         mm_interconnect_0_line7_2_s1_write;                        // mm_interconnect_0:Line7_2_s1_write -> Line7_2:write_n
	wire  [31:0] mm_interconnect_0_line7_2_s1_writedata;                    // mm_interconnect_0:Line7_2_s1_writedata -> Line7_2:writedata
	wire         mm_interconnect_0_line7_1_s1_chipselect;                   // mm_interconnect_0:Line7_1_s1_chipselect -> Line7_1:chipselect
	wire  [31:0] mm_interconnect_0_line7_1_s1_readdata;                     // Line7_1:readdata -> mm_interconnect_0:Line7_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line7_1_s1_address;                      // mm_interconnect_0:Line7_1_s1_address -> Line7_1:address
	wire         mm_interconnect_0_line7_1_s1_write;                        // mm_interconnect_0:Line7_1_s1_write -> Line7_1:write_n
	wire  [31:0] mm_interconnect_0_line7_1_s1_writedata;                    // mm_interconnect_0:Line7_1_s1_writedata -> Line7_1:writedata
	wire         mm_interconnect_0_line2_1_s1_chipselect;                   // mm_interconnect_0:Line2_1_s1_chipselect -> Line2_1:chipselect
	wire  [31:0] mm_interconnect_0_line2_1_s1_readdata;                     // Line2_1:readdata -> mm_interconnect_0:Line2_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line2_1_s1_address;                      // mm_interconnect_0:Line2_1_s1_address -> Line2_1:address
	wire         mm_interconnect_0_line2_1_s1_write;                        // mm_interconnect_0:Line2_1_s1_write -> Line2_1:write_n
	wire  [31:0] mm_interconnect_0_line2_1_s1_writedata;                    // mm_interconnect_0:Line2_1_s1_writedata -> Line2_1:writedata
	wire         mm_interconnect_0_line2_2_s1_chipselect;                   // mm_interconnect_0:LIne2_2_s1_chipselect -> LIne2_2:chipselect
	wire  [31:0] mm_interconnect_0_line2_2_s1_readdata;                     // LIne2_2:readdata -> mm_interconnect_0:LIne2_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line2_2_s1_address;                      // mm_interconnect_0:LIne2_2_s1_address -> LIne2_2:address
	wire         mm_interconnect_0_line2_2_s1_write;                        // mm_interconnect_0:LIne2_2_s1_write -> LIne2_2:write_n
	wire  [31:0] mm_interconnect_0_line2_2_s1_writedata;                    // mm_interconnect_0:LIne2_2_s1_writedata -> LIne2_2:writedata
	wire         mm_interconnect_0_line3_1_s1_chipselect;                   // mm_interconnect_0:Line3_1_s1_chipselect -> Line3_1:chipselect
	wire  [31:0] mm_interconnect_0_line3_1_s1_readdata;                     // Line3_1:readdata -> mm_interconnect_0:Line3_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line3_1_s1_address;                      // mm_interconnect_0:Line3_1_s1_address -> Line3_1:address
	wire         mm_interconnect_0_line3_1_s1_write;                        // mm_interconnect_0:Line3_1_s1_write -> Line3_1:write_n
	wire  [31:0] mm_interconnect_0_line3_1_s1_writedata;                    // mm_interconnect_0:Line3_1_s1_writedata -> Line3_1:writedata
	wire         mm_interconnect_0_line3_2_s1_chipselect;                   // mm_interconnect_0:Line3_2_s1_chipselect -> Line3_2:chipselect
	wire  [31:0] mm_interconnect_0_line3_2_s1_readdata;                     // Line3_2:readdata -> mm_interconnect_0:Line3_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line3_2_s1_address;                      // mm_interconnect_0:Line3_2_s1_address -> Line3_2:address
	wire         mm_interconnect_0_line3_2_s1_write;                        // mm_interconnect_0:Line3_2_s1_write -> Line3_2:write_n
	wire  [31:0] mm_interconnect_0_line3_2_s1_writedata;                    // mm_interconnect_0:Line3_2_s1_writedata -> Line3_2:writedata
	wire         mm_interconnect_0_line4_1_s1_chipselect;                   // mm_interconnect_0:Line4_1_s1_chipselect -> Line4_1:chipselect
	wire  [31:0] mm_interconnect_0_line4_1_s1_readdata;                     // Line4_1:readdata -> mm_interconnect_0:Line4_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line4_1_s1_address;                      // mm_interconnect_0:Line4_1_s1_address -> Line4_1:address
	wire         mm_interconnect_0_line4_1_s1_write;                        // mm_interconnect_0:Line4_1_s1_write -> Line4_1:write_n
	wire  [31:0] mm_interconnect_0_line4_1_s1_writedata;                    // mm_interconnect_0:Line4_1_s1_writedata -> Line4_1:writedata
	wire         mm_interconnect_0_line4_2_s1_chipselect;                   // mm_interconnect_0:Line4_2_s1_chipselect -> Line4_2:chipselect
	wire  [31:0] mm_interconnect_0_line4_2_s1_readdata;                     // Line4_2:readdata -> mm_interconnect_0:Line4_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line4_2_s1_address;                      // mm_interconnect_0:Line4_2_s1_address -> Line4_2:address
	wire         mm_interconnect_0_line4_2_s1_write;                        // mm_interconnect_0:Line4_2_s1_write -> Line4_2:write_n
	wire  [31:0] mm_interconnect_0_line4_2_s1_writedata;                    // mm_interconnect_0:Line4_2_s1_writedata -> Line4_2:writedata
	wire         mm_interconnect_0_line5_1_s1_chipselect;                   // mm_interconnect_0:Line5_1_s1_chipselect -> Line5_1:chipselect
	wire  [31:0] mm_interconnect_0_line5_1_s1_readdata;                     // Line5_1:readdata -> mm_interconnect_0:Line5_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line5_1_s1_address;                      // mm_interconnect_0:Line5_1_s1_address -> Line5_1:address
	wire         mm_interconnect_0_line5_1_s1_write;                        // mm_interconnect_0:Line5_1_s1_write -> Line5_1:write_n
	wire  [31:0] mm_interconnect_0_line5_1_s1_writedata;                    // mm_interconnect_0:Line5_1_s1_writedata -> Line5_1:writedata
	wire         mm_interconnect_0_line5_2_s1_chipselect;                   // mm_interconnect_0:Line5_2_s1_chipselect -> Line5_2:chipselect
	wire  [31:0] mm_interconnect_0_line5_2_s1_readdata;                     // Line5_2:readdata -> mm_interconnect_0:Line5_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line5_2_s1_address;                      // mm_interconnect_0:Line5_2_s1_address -> Line5_2:address
	wire         mm_interconnect_0_line5_2_s1_write;                        // mm_interconnect_0:Line5_2_s1_write -> Line5_2:write_n
	wire  [31:0] mm_interconnect_0_line5_2_s1_writedata;                    // mm_interconnect_0:Line5_2_s1_writedata -> Line5_2:writedata
	wire         mm_interconnect_0_line6_1_s1_chipselect;                   // mm_interconnect_0:Line6_1_s1_chipselect -> Line6_1:chipselect
	wire  [31:0] mm_interconnect_0_line6_1_s1_readdata;                     // Line6_1:readdata -> mm_interconnect_0:Line6_1_s1_readdata
	wire   [1:0] mm_interconnect_0_line6_1_s1_address;                      // mm_interconnect_0:Line6_1_s1_address -> Line6_1:address
	wire         mm_interconnect_0_line6_1_s1_write;                        // mm_interconnect_0:Line6_1_s1_write -> Line6_1:write_n
	wire  [31:0] mm_interconnect_0_line6_1_s1_writedata;                    // mm_interconnect_0:Line6_1_s1_writedata -> Line6_1:writedata
	wire         mm_interconnect_0_line6_2_s1_chipselect;                   // mm_interconnect_0:Line6_2_s1_chipselect -> Line6_2:chipselect
	wire  [31:0] mm_interconnect_0_line6_2_s1_readdata;                     // Line6_2:readdata -> mm_interconnect_0:Line6_2_s1_readdata
	wire   [1:0] mm_interconnect_0_line6_2_s1_address;                      // mm_interconnect_0:Line6_2_s1_address -> Line6_2:address
	wire         mm_interconnect_0_line6_2_s1_write;                        // mm_interconnect_0:Line6_2_s1_write -> Line6_2:write_n
	wire  [31:0] mm_interconnect_0_line6_2_s1_writedata;                    // mm_interconnect_0:Line6_2_s1_writedata -> Line6_2:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [LIne2_2:reset_n, Line1_1:reset_n, Line1_2:reset_n, Line2_1:reset_n, Line3_1:reset_n, Line3_2:reset_n, Line4_1:reset_n, Line4_2:reset_n, Line5_1:reset_n, Line5_2:reset_n, Line6_1:reset_n, Line6_2:reset_n, Line7_1:reset_n, Line7_2:reset_n, Line8_1:reset_n, Line8_2:reset_n, altpll_0:reset, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, leds:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, sdram_controller:reset_n, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	compression_LIne2_2 line2_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line2_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line2_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line2_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line2_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line2_2_s1_readdata),   //                    .readdata
		.in_port    (line2_2_in_port),                         // external_connection.export
		.out_port   (line2_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line1_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line1_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line1_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line1_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line1_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line1_1_s1_readdata),   //                    .readdata
		.in_port    (line1_1_in_port),                         // external_connection.export
		.out_port   (line1_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line1_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line1_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line1_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line1_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line1_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line1_2_s1_readdata),   //                    .readdata
		.in_port    (line1_2_in_port),                         // external_connection.export
		.out_port   (line1_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line2_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line2_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line2_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line2_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line2_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line2_1_s1_readdata),   //                    .readdata
		.in_port    (line2_1_in_port),                         // external_connection.export
		.out_port   (line2_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line3_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line3_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line3_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line3_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line3_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line3_1_s1_readdata),   //                    .readdata
		.in_port    (line3_1_in_port),                         // external_connection.export
		.out_port   (line3_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line3_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line3_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line3_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line3_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line3_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line3_2_s1_readdata),   //                    .readdata
		.in_port    (line3_2_in_port),                         // external_connection.export
		.out_port   (line3_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line4_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line4_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line4_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line4_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line4_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line4_1_s1_readdata),   //                    .readdata
		.in_port    (line4_1_in_port),                         // external_connection.export
		.out_port   (line4_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line4_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line4_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line4_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line4_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line4_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line4_2_s1_readdata),   //                    .readdata
		.in_port    (line4_2_in_port),                         // external_connection.export
		.out_port   (line4_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line5_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line5_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line5_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line5_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line5_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line5_1_s1_readdata),   //                    .readdata
		.in_port    (line5_1_in_port),                         // external_connection.export
		.out_port   (line5_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line5_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line5_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line5_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line5_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line5_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line5_2_s1_readdata),   //                    .readdata
		.in_port    (line5_2_in_port),                         // external_connection.export
		.out_port   (line5_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line6_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line6_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line6_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line6_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line6_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line6_1_s1_readdata),   //                    .readdata
		.in_port    (line6_1_in_port),                         // external_connection.export
		.out_port   (line6_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line6_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line6_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line6_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line6_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line6_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line6_2_s1_readdata),   //                    .readdata
		.in_port    (line6_2_in_port),                         // external_connection.export
		.out_port   (line6_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line7_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line7_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line7_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line7_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line7_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line7_1_s1_readdata),   //                    .readdata
		.in_port    (line7_1_in_port),                         // external_connection.export
		.out_port   (line7_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line7_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line7_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line7_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line7_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line7_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line7_2_s1_readdata),   //                    .readdata
		.in_port    (line7_2_in_port),                         // external_connection.export
		.out_port   (line7_2_out_port)                         //                    .export
	);

	compression_LIne2_2 line8_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line8_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line8_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line8_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line8_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line8_1_s1_readdata),   //                    .readdata
		.in_port    (line8_1_in_port),                         // external_connection.export
		.out_port   (line8_1_out_port)                         //                    .export
	);

	compression_LIne2_2 line8_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_line8_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_line8_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_line8_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_line8_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_line8_2_s1_readdata),   //                    .readdata
		.in_port    (line8_2_in_port),                         // external_connection.export
		.out_port   (line8_2_out_port)                         //                    .export
	);

	compression_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_clk),                                  //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	compression_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	compression_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	compression_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_w_export)                         // external_connection.export
	);

	compression_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	compression_sdram_controller sdram_controller (
		.clk            (clk_clk),                                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	compression_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	compression_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.altpll_0_pll_slave_address              (mm_interconnect_0_altpll_0_pll_slave_address),              //              altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                (mm_interconnect_0_altpll_0_pll_slave_write),                //                                .write
		.altpll_0_pll_slave_read                 (mm_interconnect_0_altpll_0_pll_slave_read),                 //                                .read
		.altpll_0_pll_slave_readdata             (mm_interconnect_0_altpll_0_pll_slave_readdata),             //                                .readdata
		.altpll_0_pll_slave_writedata            (mm_interconnect_0_altpll_0_pll_slave_writedata),            //                                .writedata
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.leds_s1_address                         (mm_interconnect_0_leds_s1_address),                         //                         leds_s1.address
		.leds_s1_write                           (mm_interconnect_0_leds_s1_write),                           //                                .write
		.leds_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                        //                                .readdata
		.leds_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                       //                                .writedata
		.leds_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                      //                                .chipselect
		.Line1_1_s1_address                      (mm_interconnect_0_line1_1_s1_address),                      //                      Line1_1_s1.address
		.Line1_1_s1_write                        (mm_interconnect_0_line1_1_s1_write),                        //                                .write
		.Line1_1_s1_readdata                     (mm_interconnect_0_line1_1_s1_readdata),                     //                                .readdata
		.Line1_1_s1_writedata                    (mm_interconnect_0_line1_1_s1_writedata),                    //                                .writedata
		.Line1_1_s1_chipselect                   (mm_interconnect_0_line1_1_s1_chipselect),                   //                                .chipselect
		.Line1_2_s1_address                      (mm_interconnect_0_line1_2_s1_address),                      //                      Line1_2_s1.address
		.Line1_2_s1_write                        (mm_interconnect_0_line1_2_s1_write),                        //                                .write
		.Line1_2_s1_readdata                     (mm_interconnect_0_line1_2_s1_readdata),                     //                                .readdata
		.Line1_2_s1_writedata                    (mm_interconnect_0_line1_2_s1_writedata),                    //                                .writedata
		.Line1_2_s1_chipselect                   (mm_interconnect_0_line1_2_s1_chipselect),                   //                                .chipselect
		.Line2_1_s1_address                      (mm_interconnect_0_line2_1_s1_address),                      //                      Line2_1_s1.address
		.Line2_1_s1_write                        (mm_interconnect_0_line2_1_s1_write),                        //                                .write
		.Line2_1_s1_readdata                     (mm_interconnect_0_line2_1_s1_readdata),                     //                                .readdata
		.Line2_1_s1_writedata                    (mm_interconnect_0_line2_1_s1_writedata),                    //                                .writedata
		.Line2_1_s1_chipselect                   (mm_interconnect_0_line2_1_s1_chipselect),                   //                                .chipselect
		.LIne2_2_s1_address                      (mm_interconnect_0_line2_2_s1_address),                      //                      LIne2_2_s1.address
		.LIne2_2_s1_write                        (mm_interconnect_0_line2_2_s1_write),                        //                                .write
		.LIne2_2_s1_readdata                     (mm_interconnect_0_line2_2_s1_readdata),                     //                                .readdata
		.LIne2_2_s1_writedata                    (mm_interconnect_0_line2_2_s1_writedata),                    //                                .writedata
		.LIne2_2_s1_chipselect                   (mm_interconnect_0_line2_2_s1_chipselect),                   //                                .chipselect
		.Line3_1_s1_address                      (mm_interconnect_0_line3_1_s1_address),                      //                      Line3_1_s1.address
		.Line3_1_s1_write                        (mm_interconnect_0_line3_1_s1_write),                        //                                .write
		.Line3_1_s1_readdata                     (mm_interconnect_0_line3_1_s1_readdata),                     //                                .readdata
		.Line3_1_s1_writedata                    (mm_interconnect_0_line3_1_s1_writedata),                    //                                .writedata
		.Line3_1_s1_chipselect                   (mm_interconnect_0_line3_1_s1_chipselect),                   //                                .chipselect
		.Line3_2_s1_address                      (mm_interconnect_0_line3_2_s1_address),                      //                      Line3_2_s1.address
		.Line3_2_s1_write                        (mm_interconnect_0_line3_2_s1_write),                        //                                .write
		.Line3_2_s1_readdata                     (mm_interconnect_0_line3_2_s1_readdata),                     //                                .readdata
		.Line3_2_s1_writedata                    (mm_interconnect_0_line3_2_s1_writedata),                    //                                .writedata
		.Line3_2_s1_chipselect                   (mm_interconnect_0_line3_2_s1_chipselect),                   //                                .chipselect
		.Line4_1_s1_address                      (mm_interconnect_0_line4_1_s1_address),                      //                      Line4_1_s1.address
		.Line4_1_s1_write                        (mm_interconnect_0_line4_1_s1_write),                        //                                .write
		.Line4_1_s1_readdata                     (mm_interconnect_0_line4_1_s1_readdata),                     //                                .readdata
		.Line4_1_s1_writedata                    (mm_interconnect_0_line4_1_s1_writedata),                    //                                .writedata
		.Line4_1_s1_chipselect                   (mm_interconnect_0_line4_1_s1_chipselect),                   //                                .chipselect
		.Line4_2_s1_address                      (mm_interconnect_0_line4_2_s1_address),                      //                      Line4_2_s1.address
		.Line4_2_s1_write                        (mm_interconnect_0_line4_2_s1_write),                        //                                .write
		.Line4_2_s1_readdata                     (mm_interconnect_0_line4_2_s1_readdata),                     //                                .readdata
		.Line4_2_s1_writedata                    (mm_interconnect_0_line4_2_s1_writedata),                    //                                .writedata
		.Line4_2_s1_chipselect                   (mm_interconnect_0_line4_2_s1_chipselect),                   //                                .chipselect
		.Line5_1_s1_address                      (mm_interconnect_0_line5_1_s1_address),                      //                      Line5_1_s1.address
		.Line5_1_s1_write                        (mm_interconnect_0_line5_1_s1_write),                        //                                .write
		.Line5_1_s1_readdata                     (mm_interconnect_0_line5_1_s1_readdata),                     //                                .readdata
		.Line5_1_s1_writedata                    (mm_interconnect_0_line5_1_s1_writedata),                    //                                .writedata
		.Line5_1_s1_chipselect                   (mm_interconnect_0_line5_1_s1_chipselect),                   //                                .chipselect
		.Line5_2_s1_address                      (mm_interconnect_0_line5_2_s1_address),                      //                      Line5_2_s1.address
		.Line5_2_s1_write                        (mm_interconnect_0_line5_2_s1_write),                        //                                .write
		.Line5_2_s1_readdata                     (mm_interconnect_0_line5_2_s1_readdata),                     //                                .readdata
		.Line5_2_s1_writedata                    (mm_interconnect_0_line5_2_s1_writedata),                    //                                .writedata
		.Line5_2_s1_chipselect                   (mm_interconnect_0_line5_2_s1_chipselect),                   //                                .chipselect
		.Line6_1_s1_address                      (mm_interconnect_0_line6_1_s1_address),                      //                      Line6_1_s1.address
		.Line6_1_s1_write                        (mm_interconnect_0_line6_1_s1_write),                        //                                .write
		.Line6_1_s1_readdata                     (mm_interconnect_0_line6_1_s1_readdata),                     //                                .readdata
		.Line6_1_s1_writedata                    (mm_interconnect_0_line6_1_s1_writedata),                    //                                .writedata
		.Line6_1_s1_chipselect                   (mm_interconnect_0_line6_1_s1_chipselect),                   //                                .chipselect
		.Line6_2_s1_address                      (mm_interconnect_0_line6_2_s1_address),                      //                      Line6_2_s1.address
		.Line6_2_s1_write                        (mm_interconnect_0_line6_2_s1_write),                        //                                .write
		.Line6_2_s1_readdata                     (mm_interconnect_0_line6_2_s1_readdata),                     //                                .readdata
		.Line6_2_s1_writedata                    (mm_interconnect_0_line6_2_s1_writedata),                    //                                .writedata
		.Line6_2_s1_chipselect                   (mm_interconnect_0_line6_2_s1_chipselect),                   //                                .chipselect
		.Line7_1_s1_address                      (mm_interconnect_0_line7_1_s1_address),                      //                      Line7_1_s1.address
		.Line7_1_s1_write                        (mm_interconnect_0_line7_1_s1_write),                        //                                .write
		.Line7_1_s1_readdata                     (mm_interconnect_0_line7_1_s1_readdata),                     //                                .readdata
		.Line7_1_s1_writedata                    (mm_interconnect_0_line7_1_s1_writedata),                    //                                .writedata
		.Line7_1_s1_chipselect                   (mm_interconnect_0_line7_1_s1_chipselect),                   //                                .chipselect
		.Line7_2_s1_address                      (mm_interconnect_0_line7_2_s1_address),                      //                      Line7_2_s1.address
		.Line7_2_s1_write                        (mm_interconnect_0_line7_2_s1_write),                        //                                .write
		.Line7_2_s1_readdata                     (mm_interconnect_0_line7_2_s1_readdata),                     //                                .readdata
		.Line7_2_s1_writedata                    (mm_interconnect_0_line7_2_s1_writedata),                    //                                .writedata
		.Line7_2_s1_chipselect                   (mm_interconnect_0_line7_2_s1_chipselect),                   //                                .chipselect
		.Line8_1_s1_address                      (mm_interconnect_0_line8_1_s1_address),                      //                      Line8_1_s1.address
		.Line8_1_s1_write                        (mm_interconnect_0_line8_1_s1_write),                        //                                .write
		.Line8_1_s1_readdata                     (mm_interconnect_0_line8_1_s1_readdata),                     //                                .readdata
		.Line8_1_s1_writedata                    (mm_interconnect_0_line8_1_s1_writedata),                    //                                .writedata
		.Line8_1_s1_chipselect                   (mm_interconnect_0_line8_1_s1_chipselect),                   //                                .chipselect
		.Line8_2_s1_address                      (mm_interconnect_0_line8_2_s1_address),                      //                      Line8_2_s1.address
		.Line8_2_s1_write                        (mm_interconnect_0_line8_2_s1_write),                        //                                .write
		.Line8_2_s1_readdata                     (mm_interconnect_0_line8_2_s1_readdata),                     //                                .readdata
		.Line8_2_s1_writedata                    (mm_interconnect_0_line8_2_s1_writedata),                    //                                .writedata
		.Line8_2_s1_chipselect                   (mm_interconnect_0_line8_2_s1_chipselect),                   //                                .chipselect
		.onchip_memory2_0_s1_address             (mm_interconnect_0_onchip_memory2_0_s1_address),             //             onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write               (mm_interconnect_0_onchip_memory2_0_s1_write),               //                                .write
		.onchip_memory2_0_s1_readdata            (mm_interconnect_0_onchip_memory2_0_s1_readdata),            //                                .readdata
		.onchip_memory2_0_s1_writedata           (mm_interconnect_0_onchip_memory2_0_s1_writedata),           //                                .writedata
		.onchip_memory2_0_s1_byteenable          (mm_interconnect_0_onchip_memory2_0_s1_byteenable),          //                                .byteenable
		.onchip_memory2_0_s1_chipselect          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),          //                                .chipselect
		.onchip_memory2_0_s1_clken               (mm_interconnect_0_onchip_memory2_0_s1_clken),               //                                .clken
		.sdram_controller_s1_address             (mm_interconnect_0_sdram_controller_s1_address),             //             sdram_controller_s1.address
		.sdram_controller_s1_write               (mm_interconnect_0_sdram_controller_s1_write),               //                                .write
		.sdram_controller_s1_read                (mm_interconnect_0_sdram_controller_s1_read),                //                                .read
		.sdram_controller_s1_readdata            (mm_interconnect_0_sdram_controller_s1_readdata),            //                                .readdata
		.sdram_controller_s1_writedata           (mm_interconnect_0_sdram_controller_s1_writedata),           //                                .writedata
		.sdram_controller_s1_byteenable          (mm_interconnect_0_sdram_controller_s1_byteenable),          //                                .byteenable
		.sdram_controller_s1_readdatavalid       (mm_interconnect_0_sdram_controller_s1_readdatavalid),       //                                .readdatavalid
		.sdram_controller_s1_waitrequest         (mm_interconnect_0_sdram_controller_s1_waitrequest),         //                                .waitrequest
		.sdram_controller_s1_chipselect          (mm_interconnect_0_sdram_controller_s1_chipselect),          //                                .chipselect
		.sysid_qsys_control_slave_address        (mm_interconnect_0_sysid_qsys_control_slave_address),        //        sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata       (mm_interconnect_0_sysid_qsys_control_slave_readdata)        //                                .readdata
	);

	compression_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
